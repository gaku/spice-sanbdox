* Zener Diode Voltage Regulator
Vin 1 0 DC 9V
R1 1 2 47
* 'zener' is a model name
D1 0 2 zener
* Model definition of 'zener' diode. BV is reverse breakdown voltage.
.model zener D (BV=3.3V)
.control
** DC from 0V to 9V with 0.5V increment
dc Vin 0 5 0.1
print v(1) i(Vin) v(2)
.endc
.end
